`timescale 1ns/10ps

`ifdef syn
`include "/usr/cad/CBDK/Executable_Package/Collaterals/IP/stdcell/N16ADFP_StdCell/VERILOG/N16ADFP_StdCell.v"
`include "ALU_syn.v"
`else
`include "ALU.v"
`endif

`define DATA_SIZE  32
`define OP_SIZE  5

`define ADD    5'b00000
`define SUB    5'b00001
`define OR     5'b00010
`define AND    5'b00011
`define XOR    5'b00100
`define NOT    5'b00101
`define NAND   5'b00110
`define NOR    5'b00111
`define SLT    5'b01000
`define SLTU   5'b01001
`define ABS    5'b01010
`define BITREV 5'b01011

module tb_ALU;

// ----------------------   reg   ---------------------- //
reg   [`OP_SIZE-1:0]  alu_op1;
reg   [`DATA_SIZE-1:0]   src1;
reg   [`DATA_SIZE-1:0]   src2;

// ----------------------   wire  ---------------------- //
wire   [`DATA_SIZE-1:0]  alu_out1;
wire                    alu_overflow1;

integer error;
integer i;

ALU ALU (
	.alu_op(alu_op1),
	.src1(src1),
	.src2(src2),
    .alu_out(alu_out1),
	.alu_overflow(alu_overflow1)
);

initial begin
	$monitor($time, " opcode1 = %h, src1 = %h, src2 = %h, alu_out = %h, alu_overflow = %h ", alu_op1,  src1, src2, alu_out1, alu_overflow1);
end

initial begin
	error=0;
	#5
	if(alu_out1==32'h0000_0011 && alu_overflow1==1'b0 )begin//ADD1
		error = error;
	end
	else begin
		$display("there are some errors with ADD ");
		$finish;
		error = error +1;
	end
	#10
	if(alu_out1==32'h0000_0001 && alu_overflow1==1'b0 )begin//ADD2
		error = error;
	end
	else begin
		$display("there are some errors with ADD  ");
		$finish;
		error = error +1;
	end
	#10
	if(alu_out1==32'h8000_0001 && alu_overflow1==1'b1 ) begin//ADD3
		error = error;
	end
	else begin
		$display("there are some errors with ADD  ");
		$finish;
		error = error +1;
	end
	#10
	if(alu_out1==32'hffff_ffff && alu_overflow1==1'b0  )begin//SUB
		error = error;
	end
	else begin
		$display("there are some errors with SUB ");
		$finish;
		error = error +1;
	end
	#10
	if(alu_out1==32'hffff_0000 && alu_overflow1==1'b0 )begin //OR
		error = error;
	end
	else begin
		$display("there are some errors with OR  ");
		$finish;
		error = error +1;
	end
	#10
	if(alu_out1==32'h00ff_0000 && alu_overflow1==1'b0 )begin//AND 
		error = error;
	end
	else begin
		
		$display("there are some errors with AND  ");
		$finish;
		error = error +1;
	end
	#10
	if(alu_out1==32'hff00_ff00 && alu_overflow1==1'b0 )begin//XOR 
		error = error;
	end
	else begin
		$display("there are some errors with XOR");
		$finish;
		error = error +1;
	end
	#10
	if(alu_out1==32'hffff_0000 && alu_overflow1==1'b0)begin//NOT
		error = error;
	end
	else begin
		
		$display("there are some errors with NOT ");
		$finish;
		error = error +1;
	end
	#10
	if(alu_out1==32'hff00_ffff && alu_overflow1==1'b0 )begin//NAND 
		error = error;
	end
	else begin
		$display("there are some errors with NAND");
		$finish;
		error = error +1;
	end
	#10
	if(alu_out1==32'h0000_ffff && alu_overflow1==1'b0)begin//NOR
		error = error;
	end
	else begin
		
		$display("there are some errors with NOR ");
		$finish;
		error = error +1;
	end
	
	//---------------------------------------------------------
	#10
	if(alu_out1==32'h0000_0000 && alu_overflow1==1'b0 )begin//SLT
		error = error;
	end
	else begin
		$display("there are some errors with SLT");
		$finish;
		error = error +1;
	end
	#10
	if(alu_out1==32'h0000_0001 && alu_overflow1==1'b0 )begin//SLTU
		error = error;
	end
	else begin
		$display("there are some errors with SLTU");
		$finish;
		error = error +1;
	end
	#10
	if(alu_out1==32'h0000_0087 && alu_overflow1==1'b0 )begin//ABS
		error = error;
	end
	else begin
		$display("there are some errors with ABS");
		$finish;
		error = error +1;
	end
	#10
	if(alu_out1==32'h0000_0003 && alu_overflow1==1'b0 )begin//BITREV 
		error = error;
	end
	else begin
		$display("there are some errors with BITREV ");
		$finish;
		error = error +1;
	end
	#10
  
	if(error === 0)begin
		$display("\n");
        $display("\n");
for(i=0;i<=5000;i=i+1) begin
	if(i%2==0) begin
$display("	     ,(((((((((())))))))),	      ");
$display("	   ,((((((((((()))))))))))),	      ");
$display("	  ,(((((((((\\\|///))))))))),	      ");
$display("	 ,((((((((((///|\\\)))))))))),	  ");
$display("	 ((((((((//////^\\\\\\))))))))	  ");
$display("	 ((((((' .-\"\"-   -\"\"-. '))))))  ");
$display("	 (((((  `\.-.     .-./`  )))))	  ");
$display("	 ((((( -=(0) )   (0) )=- )))))	  ");
$display("	 '((((   /'-'     '-'\\   ))))'	  ");
$display("	  ((((\   _,   A  ,_    /))))	      ");
$display("	  '((((\    \     /    /))))'	      ");
$display("	    '((('.   `-o-'   .')))'	      ");
$display("	          '-.,___,.-'				  ");
	end
	else begin
$display("					     ,(((((((((())))))))),	      ");
$display("					   ,((((((((((()))))))))))),	      ");
$display("					  ,(((((((((\\\|///))))))))),	      ");
$display("					 ,((((((((((///|\\\)))))))))),	  ");
$display("					 ((((((((//////^\\\\\\))))))))	  ");
$display("					 ((((((' .-\"\"-   -\"\"-. '))))))  ");
$display("					 (((((  `\.-.     .-./`  )))))	  ");
$display("					 ((((( -=(0) )   (0) )=- )))))	  ");
$display("					 '((((   /'-'     '-'\\   ))))'	  ");
$display("					  ((((\   _,   A  ,_    /))))	      ");
$display("					  '((((\    \     /    /))))'	      ");
$display("					    '((('.   `-o-'   .')))'	      ");
$display("					          '-.,___,.-'				  ");		
	end
end

$display("					     ,(((((((((())))))))),	      ");
$display("					   ,((((((((((()))))))))))),	      ");
$display("					  ,(((((((((\\\|///))))))))),	      ");
$display("					 ,((((((((((///|\\\)))))))))),	  ");
$display("					 ((((((((//////^\\\\\\))))))))	  ");
$display("					 ((((((' .-\"\"-   -\"\"-. '))))))  ");
$display("					 (((((  `\.-.     .-./`  )))))	  ");
$display("					 ((((( -=(0) )   (0) )=- )))))	  ");
$display("					 '((((   /'-'     '-'\\   ))))'	  ");
$display("					  ((((\   _,   A  ,_    /))))	      ");
$display("					  '((((\    \     /    /))))'	      ");
$display("					    '((('.   `-o-'   .')))'	      ");
$display("					          '-.,___,.-'				  ");
$display("\n");
$display(" ppppp   ppppppppp     aaaaaaaaaaaaa      ssssssssss       ssssssssss   ");
$display(" p::::ppp:::::::::p    a::::::::::::a   ss::::::::::s    ss::::::::::s  ");
$display(" p:::::::::::::::::p   aaaaaaaaa:::::ass:::::::::::::s ss:::::::::::::s ");
$display(" pp::::::ppppp::::::p           a::::as::::::ssss:::::ss::::::ssss:::::s");
$display("  p:::::p     p:::::p    aaaaaaa:::::a s:::::s  ssssss  s:::::s  ssssss ");
$display("  p:::::p     p:::::p  aa::::::::::::a   s::::::s         s::::::s      ");
$display("  p:::::p     p:::::p a::::aaaa::::::a      s::::::s         s::::::s   ");
$display("  p:::::p    p::::::pa::::a    a:::::assssss   s:::::s ssssss   s:::::s ");
$display("  p:::::ppppp:::::::pa::::a    a:::::as:::::ssss::::::ss:::::ssss::::::s");
$display("  p::::::::::::::::p a:::::aaaa::::::as::::::::::::::s s::::::::::::::s ");
$display("  p::::::::::::::pp   a::::::::::aa:::as:::::::::::ss   s:::::::::::ss  ");
$display("  p::::::pppppppp      aaaaaaaaaa  aaaa sssssssssss      sssssssssss    ");
$display("  p:::::p                                                               ");
$display("  p:::::p                                                               ");
$display(" ppppppppp                                                              ");
$display("	     ,(((((((((())))))))),	      ");
$display("	   ,((((((((((()))))))))))),	      ");
$display("	  ,(((((((((\\\|///))))))))),	      ");
$display("	 ,((((((((((///|\\\)))))))))),	  ");
$display("	 ((((((((//////^\\\\\\))))))))	  ");
$display("	 ((((((' .-\"\"-   -\"\"-. '))))))  ");
$display("	 (((((  `\.-.     .-./`  )))))	  ");
$display("	 ((((( -=(0) )   (0) )=- )))))	  ");
$display("	 '((((   /'-'     '-'\\   ))))'	  ");
$display("	  ((((\   _,   A  ,_    /))))	      ");
$display("	  '((((\    \     /    /))))'	      ");
$display("	    '((('.   `-o-'   .')))'	      ");
$display("	          '-.,___,.-'				  ");
$display("\n");
	end
	else begin
$display("\n");
$display("\n");
$display("			  `-.     `.   \      :      /   .'     .-'					");
$display("			     `-.    `.  `.    :    .'  .'    .-'   				");
$display("			 `-._   `-.   `.  \   :   /  .'   .-'   _.-		");
$display("			 _   `-._  `-.  `. `. : .' .'  .-'  _.-'   				");
$display("			  `--._  `-._ `-. `. \:/ .' .-' _.-'  _.--'				");
$display("			 .__   `--._ `-._`-.`_=_'.-'_.-' _.--'   __			");
$display("			 _  `--.__  `--._`-q(-_-)p-'_.--'  __.--'  				");
$display("			  `--..__ `--.__ `-'_) (_`-' __.--' __..--'		");
$display("			 `--..__ `--..__`--/__/  \--'__..--' __..--				");
$display("			 ___    ``--..__`_(<_   _/)_'__..--''    __		");
$display("			 ___```---...___(__\_\_|_/__)___...---'''__				");
$display("\n");
$display("                              OOPS! Simulation Failed !!");
$display("\n");
$display("\n");
    end
end

initial begin
	#0	alu_op1 = `ADD;  	src1 = 32'h0000_000f; src2 = 32'h0000_0002;// 15 , 2, 0000_0011
	#10	alu_op1 = `ADD;  	src1 = 32'hffff_ffff; src2 = 32'h0000_0002;// -1 , 2, 0000_0001,ffff_fffd
	#10	alu_op1 = `ADD;  	src1 = 32'h7fff_ffff; src2 = 32'h0000_0002;// overflow, 8000_0001 ,ffff_fffe
	#10	alu_op1 = `SUB;  	src1 = 32'h0000_0001; src2 = 32'h0000_0002;// 1 , 2, ffff_ffff,0000_0003
	#10	alu_op1 = `OR;		src1 = 32'hffff_0000; src2 = 32'h0000_0000;// ffff_0000 ,0000_0000
	#10	alu_op1 = `AND;  	src1 = 32'hffff_0000; src2 = 32'h00ff_0000;// 00ff_0000 ,00fe_0000
	#10	alu_op1 = `XOR;  	src1 = 32'hffff_0000; src2 = 32'h00ff_ff00;// ff00_ff00 ,ff00_ff00
	#10 alu_op1 = `NOT;  	src1 = 32'h0000_ffff; src2 = 32'h0000_0000;// ffff_0000 ,0000_ffff
	#10 alu_op1 = `NAND; 	src1 = 32'hffff_0000; src2 = 32'h00ff_0000;// ff00_ffff ,ff00_ffff
	#10 alu_op1 = `NOR;  	src1 = 32'hffff_0000; src2 = 32'h0000_0000;// 0000_ffff ,0000_ffff
	#10	alu_op1 = `SLT;  	src1 = 32'h1234_5678; src2 = 32'hffff_ffff;// 0000_0000 ,0000_0000
	#10	alu_op1 = `SLTU; 	src1 = 32'h1234_5678; src2 = 32'hffff_ffff;// 0000_0001 ,0000_0001
	#10 alu_op1 = `ABS;  	src1 = 32'hffff_ff79; src2 = 32'h0000_0000;// |-135| = 135
	#10 alu_op1 = `BITREV;  src1 = 32'hc000_0000; src2 = 32'h0000_0000;// 0000_0003, 3fff_ffff
	
	#100  $finish;
end

initial begin
	`ifdef FSDB
		$fsdbDumpfile("ALU.fsdb");
		$fsdbDumpvars;
	`endif
end

`ifdef syn
	initial $sdf_annotate("ALU_syn.sdf", ALU);
`endif

endmodule
