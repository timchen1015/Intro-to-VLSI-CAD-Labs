module HA (
    input a ,
    input b ,
    output sum ,
    output carry
);

//put your design here
    
endmodule